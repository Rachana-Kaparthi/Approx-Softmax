module LOD32 ( input [31:0] data,
                output [4:0] sel);

assign sel[4] = (data[31:16]==0) ? 0:1;
assign sel[3] = (sel[4]) ? ((data[31:24]==0) ? 0:1) : ((data[15:8]==0) ? 0:1);
assign sel[2] = (sel[4]) ? ((sel[3]) ? ((data[31:28]==0) ? 0:1) : ((data[23:20]==0) ? 0:1)) : ((sel[3]) ? ((data[15:12]==0) ? 0:1) : ((data[7:4]==0) ? 0:1));
assign sel[1] = (sel[4]) ? ((sel[3]) ? ((sel[2]) ? ((data[31:30]==0) ? 0:1) : ((data[27:26]==0) ? 0:1)) : ((sel[2]) ? ((data[23:22]==0) ? 0:1) : ((data[19:18]==0) ? 0:1))) : ((sel[3]) ? ((sel[2]) ? ((data[15:14]==0) ? 0:1) : ((data[11:10]==0) ? 0:1)) : ((sel[2]) ? ((data[7:6]==0) ? 0:1) : ((data[3:2]==0) ? 0:1)));
assign sel[0] = (sel[4]) ? ((sel[3]) ? ((sel[2]) ? ((sel[1]) ? ((data[31]==0) ? 0:1) : ((data[29]==0) ? 0:1)) : ((sel[1]) ? ((data[27]==0) ? 0:1) : ((data[25]==0) ? 0:1))) : ((sel[2]) ? ((sel[1]) ? ((data[23]==0) ? 0:1) : ((data[21]==0) ? 0:1)) : ((sel[1]) ? ((data[19]==0) ? 0:1) : ((data[17]==0) ? 0:1)))) : ((sel[3]) ? ((sel[2]) ? ((sel[1]) ? ((data[15]==0) ? 0:1) : ((data[13]==0) ? 0:1)) : ((sel[1]) ? ((data[11]==0) ? 0:1) : ((data[9]==0) ? 0:1))) : ((sel[3]) ? ((sel[2]) ? ((data[7]==0) ? 0:1) : ((data[5]==0) ? 0:1)) : ((sel[1]) ? ((data[3]==0) ? 0:1) : ((data[1]==0) ? 0:1))));

endmodule




module LOD64(
output [5:0] sel,
input [63:0]data );


assign sel[5] =  (data[63:32] == 0) ? 0 :1;
assign sel[4] = (sel[5] ) ? ((data[63:48] == 0) ? 0 : 1) : ((data[31:16] == 0) ? 0:1);
assign sel[3] = (sel[5]) ? ((sel[4]) ? ((data[63:56] ==0) ? 0:1) : ((data[47:40]==0) ? 0:1)) : ((sel[4]) ? ((data[31:24] ==0) ? 0:1) : ((data[15:8]==0) ? 0:1));
assign sel[2] = (sel[5]) ? ((sel[4]) ? ((sel[3]) ? ((data[63:60] == 0) ? 0:1) : ((data[55:52] ==0)? 0:1)) : ((sel[3]) ? ((data[47:44] == 0 ? 0:1)) : ((data[39:36] == 0 ?0:1)))) : ((sel[4]) ? ((sel[3]) ? ((data[31:28] == 0) ? 0:1) : ((data[23:20] ==0)? 0:1)) : ((sel[3]) ? ((data[15:12] == 0 ? 0:1)) : ((data[7:4] == 0 ?0:1))));
//assign sel[1] = (sel[5]) ? ((sel[4]) ? ((sel[3]) ? (((sel[2]) ? ((data[63:62]==0) ? 0:1) : ((data[59:58]==0) ? 0:1)) : ((sel[2]) ? ((data[55:54]==0) ? 0:1) : ((data[51:50]==0) ? 0:1))) : ((sel[3]) ? (((sel[2]) ? ((data[47:46]==0) ? 0:1) : ((data[43:42]==0) ? 0:1)) : ((sel[2]) ? ((data[39:38]==0) ? 0:1) : ((data[35:34]==0) ? 0:1))) ))) : ((sel[4]) ? ((sel[3]) ? (((sel[2]) ? ((data[31:30]==0) ? 0:1) : ((data[27:26]==0) ? 0:1)) : ((sel[2]) ? ((data[23:22]==0) ? 0:1) : ((data[19:18]==0) ? 0:1))) : ((sel[3]) ? (((sel[2]) ? ((data[15:14]==0) ? 0:1) : ((data[11:10]==0) ? 0:1)) : ((sel[2]) ? ((data[7:6]==0) ? 0:1) : ((data[3:2]==0) ? 0:1))) )));
//assign sel[0] = (sel[5] ? ((sel[4]) ? ((sel[3]) ? ((sel[2]) ? ((sel[1]) ? ((data[63]==0) ? 0:1) : ((data[61]==0) ? 0:1)) : ((sel[1]) ? ((data[59]==0) ? 0:1) : ((data[57]==0) ? 0:1))) : ((sel[2]) ? ((sel[1]) ? ((data[55]==0) ? 0:1) : ((data[53]==0) ? 0:1)) : ((sel[1]) ? ((data[51]==0) ? 0:1) : ((data[49]==0) ? 0:1))) : ((sel[3]) ? ((sel[2]) ? ((sel[1]) ? ((data[47]==0) ? 0:1) : ((data[45]==0) ? 0:1)) : ((sel[1]) ? ((data[43]==0) ? 0:1) : ((data[41]==0) ? 0:1))) : ((sel[2]) ? ((sel[1]) ? ((data[39]==0) ? 0:1) : ((data[37]==0) ? 0:1)) : ((sel[1]) ? ((data[35]==0) ? 0:1) : ((data[33]==0) ? 0:1))) : ((sel[4]) ? ((sel[3]) ? ((sel[2]) ? ((sel[1]) ? ((data[31]==0) ? 0:1) : ((data[29]==0) ? 0:1)) : ((sel[1]) ? ((data[27]==0) ? 0:1) : ((data[25]==0) ? 0:1))) : ((sel[2]) ? ((sel[1]) ? ((data[23]==0) ? 0:1) : ((data[21]==0) ? 0:1)) : ((sel[1]) ? ((data[19]==0) ? 0:1) : ((data[17]==0) ? 0:1))) : ((sel[3]) ? ((sel[2]) ? ((sel[1]) ? ((data[15]==0) ? 0:1) : ((data[13]==0) ? 0:1)) : ((sel[1]) ? ((data[11]==0) ? 0:1) : ((data[9]==0) ? 0:1))) : ((sel[2]) ? ((sel[1]) ? ((data[7]==0) ? 0:1) : ((data[5]==0) ? 0:1)) : ((sel[1]) ? ((data[3]==0) ? 0:1) : ((data[1]==0) ? 0:1))) )) )))));
assign sel[1] = (sel[5]) ? ((sel[4]) ? ((sel[3]) ? ((sel[2]) ? ((data[63:62]==0) ? 0:1) : ((data[59:58]==0) ? 0:1)) : ((sel[2]) ? ((data[55:54]==0) ? 0:1) : ((data[51:50]==0) ? 0:1)) ):((sel[3]) ? ((sel[2]) ? ((data[47:46]==0) ? 0:1) : ((data[43:42]==0) ? 0:1)) : ((sel[2]) ? ((data[39:38]==0) ? 0:1) : ((data[35:34]==0) ? 0:1)) )) : ((sel[4]) ? ((sel[3]) ? ((sel[2]) ? ((data[31:30]==0) ? 0:1): ((data[27:26]==0) ? 0:1)) : ((sel[2]) ? ((data[23:22]==0) ? 0:1) : ((data[19:18]==0) ? 0:1))) : ((sel[3]) ? ((sel[2]) ? ((data[15:14]==0) ? 0:1) : ((data[11:10]==0) ? 0:1)) : ((sel[2]) ? ((data[7:6]==0) ? 0:1) : ((data[3:2]==0) ? 0:1))) ); 
assign sel[0] = (sel[5]) ?  
                ((sel[4]) ? ((sel[3]) ? ((sel[2]) ? ((sel[1]) ? ((data[63]==0) ? 0:1) : ((data[61]==0) ? 0:1)) : ((sel[1]) ? ((data[59]==0) ? 0:1) : ((data[57]==0) ? 0:1))) : ((sel[2]) ? ((sel[1]) ? ((data[55]==0) ? 0:1) : ((data[53]==0) ? 0:1)) : ((sel[1]) ? ((data[51]==0) ? 0:1) : ((data[49]==0) ? 0:1)))) : ((sel[3]) ? ((sel[2]) ? ((sel[1]) ? ((data[47]==0) ? 0:1) : ((data[45]==0) ? 0:1)) : ((sel[1]) ? ((data[43]==0) ? 0:1) : ((data[41]==0) ? 0:1))) : ((sel[2]) ? ((sel[1]) ? ((data[39]==0) ? 0:1) : ((data[37]==0) ? 0:1)) : ((sel[1]) ? ((data[35]==0) ? 0:1): ((data[33]==0) ? 0:1))))):
                ((sel[4]) ? ((sel[3]) ? ((sel[2]) ? ((sel[1]) ? ((data[31]==0) ? 0:1) : ((data[29]==0) ? 0:1)) : ((sel[1]) ? ((data[27]==0) ? 0:1) : ((data[25]==0) ? 0:1))) : ((sel[2]) ? ((sel[1]) ? ((data[23]==0) ? 0:1) : ((data[21]==0) ? 0:1)) : ((sel[1]) ? ((data[19]==0) ? 0:1) : ((data[17]==0) ? 0:1)))) : ((sel[3]) ? ((sel[2]) ? ((sel[1]) ? ((data[15]==0) ? 0:1) : ((data[13]==0) ? 0:1)) : ((sel[1]) ? ((data[11]==0) ? 0:1) : ((data[9] ==0) ? 0:1))) : ((sel[2]) ? ((sel[1]) ? ((data[7]==0) ? 0:1) : ((data[5]==0) ? 0:1)) : ((sel[1]) ? ((data[3]==0) ? 0:1) : ((data[1]==0) ? 0:1)))));

endmodule
